library verilog;
use verilog.vl_types.all;
entity Lab6_testbench is
end Lab6_testbench;
