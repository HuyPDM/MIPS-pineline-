library verilog;
use verilog.vl_types.all;
entity Counter_testbench is
end Counter_testbench;
